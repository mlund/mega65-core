use WORK.ALL;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use Std.TextIO.all;
use work.debugtools.all;
use work.cputypes.all;

-- on Pi1541 test unit:
-- ATN - purple
-- SRQ - white
-- DATA - green
-- CLK - blue

entity iec_serial is
  generic (
    cpu_frequency : integer
    );
  port (
    clock : in std_logic;
    clock81 : in std_logic;
    irq : out std_logic := '1';
    
    --------------------------------------------------
    -- CBM floppy serial port
    --------------------------------------------------
    fastio_addr : in unsigned(19 downto 0);
    fastio_write : in std_logic;
    fastio_read : in std_logic;
    fastio_wdata : in unsigned(7 downto 0);
    fastio_rdata : out unsigned(7 downto 0);

    debug_state : out unsigned(11 downto 0);
    debug_usec : out unsigned(7 downto 0);
    debug_msec : out unsigned(7 downto 0);
    debug_waits : out unsigned(7 downto 0);
    iec_state_reached : out unsigned(11 downto 0);
    
    --------------------------------------------------
    -- CBM floppy serial port
    --------------------------------------------------
    iec_reset : out std_logic := '1';
    iec_atn : out std_logic;
    iec_clk_en : out std_logic;
    iec_data_en : out std_logic;
    iec_srq_en : out std_logic;
    iec_clk_o : out std_logic;
    iec_data_o : out std_logic;
    iec_srq_o : out std_logic;
    iec_clk_i : in std_logic;
    iec_data_i : in std_logic;
    iec_srq_i : in std_logic
    
    );
end iec_serial;

architecture questionable of iec_serial is

  signal iec_irq : unsigned(7 downto 0) := x"00";
  signal iec_status : unsigned(7 downto 0) := x"00";
  signal iec_data : unsigned(7 downto 0) := x"00";
  signal iec_data_out : unsigned(7 downto 0) := x"00";
  signal iec_devinfo : unsigned(7 downto 0) := x"00";

  signal iec_cmd : unsigned(7 downto 0) := x"00";
  signal iec_new_cmd : std_logic := '0';

  -- C= fast serial protocol does not send fast byte prior
  -- to ATN if a device is listening (as in that case, it
  -- would treat the byte as data)
  signal iec_dev_listening : std_logic := '0';  
  
  signal iec_state : integer := 0;
  signal last_iec_state : integer := 0;
  signal iec_busy : std_logic := '0';
  signal iec_under_attention : std_logic := '0';
  
  signal wait_clk_high : std_logic := '0';
  signal wait_clk_low : std_logic := '0';
  signal wait_data_high : std_logic := '0';
  signal wait_data_low : std_logic := '0';
  signal wait_srq_high : std_logic := '0';
  signal wait_srq_low : std_logic := '0';

  signal wait_usec : integer := 0;
  signal wait_msec : integer := 0;

  signal iec_advance : std_logic := '0';

  signal cycles : integer := 0;
  signal usecs : integer := 0;
  signal usec_toggle : std_logic := '0';
  signal msec_toggle : std_logic := '0';
  signal last_usec_toggle : std_logic := '0';
  signal last_msec_toggle : std_logic := '0';
  signal timing_sync_toggle : std_logic := '0';
  signal last_timing_sync_toggle : std_logic := '0';

  signal last_iec_data : std_logic := 'U';
  signal last_iec_clk : std_logic := 'U';
  signal last_iec_srq : std_logic := 'U';
  
begin

  -- Note that we put RX on bit 6, so that the common case of LOADing can be a
  -- little faster, by allowing BIT $D697 / BVC *-3 to be a very tight loop
  -- for waiting for bytes.

  -- @IO:GS $D697.7 AUTOIEC:IRQFLAG Interrupt flag. Set if any IRQ event is triggered.
  -- @IO:GS $D697.6 AUTOIEC:IRQRX Set if a byte has been received from a listener.
  -- @IO:GS $D697.5 AUTOIEC:IRQREADY Set if ready to process a command
  -- @IO:GS $D697.4 AUTOIEC:IRQTO Set if a protocol timeout has occurred, e.g., device not found.
  -- @IO:GS $D697.3 AUTOIEC:IRQEN Enable interrupts if set
  -- @IO:GS $D697.2 AUTOIEC:IRQRXEN Enable RX interrupt source if set
  -- @IO:GS $D697.1 AUTOIEC:IRQREADYEN Enable TX interrupt source if set
  -- @IO:GS $D697.0 AUTOIEC:IRQTOEN Enable timeout interrupt source if set
  
  -- @IO:GS $D698.7 AUTOIEC:STNODEV Device not present
  -- @IO:GS $D698.6 AUTOIEC:STNOEOF End of file
  -- @IO:GS $D698.5 AUTOIEC:STSRQ State of SRQ line
  -- @IO:GS $D698.4 AUTOIEC:STVERIFY Verify error occurred
  -- @IO:GS $D698.3 AUTOIEC:STC State of CLK line
  -- @IO:GS $D698.2 AUTOIEC:STD Sate of DATA line
  -- @IO:GS $D698.1 AUTOIEC:STTO Timeout occurred
  -- @IO:GS $D698.0 AUTOIEC:STDDIR Data direction when timeout occurred.
  
  -- @IO:GS $D699 AUTOIEC:DATA Data byte read from IEC bus
  -- @IO:GS $D69A.7 AUTOIEC:DIPRESENT Device is present
  -- @IO:GS $D69A.5-6 AUTOIEC:DIPROT Device protocol (00=1541,01=C128/C65 FAST, 10 = JiffyDOS(tm), 11=both
  -- @IO:GS $D69A.4 AUTOIEC:DIATN Device is currently held under attention
  -- @IO:GS $D69A.0-3 AUTOIEC:DIDEVNUM Lower 4 bits of currently selected device number
  
  process (clock,clock81) is
    procedure d(v : std_logic) is
    begin
      if v /= last_iec_data then
        report "SIGNAL: Setting DATA to " & std_logic'image(v);
        last_iec_data <= v;
      end if;
      iec_data_o <= v; iec_data_en <= v;      
    end procedure;
    procedure c(v : std_logic) is
    begin
      if v /= last_iec_clk then
        report "SIGNAL: Setting CLK to " & std_logic'image(v);
        last_iec_clk <= v;
      end if;
      iec_clk_o <= v; iec_clk_en <= v;      
    end procedure;
    procedure s(v : std_logic) is
    begin
      if v/= last_iec_srq then
        report "SIGNAL: Setting SRQ to " & std_logic'image(v);
        last_iec_srq <= v;
      end if;
      iec_srq_o <= v; iec_srq_en <= v;      
    end procedure;
    procedure a(v : std_logic) is
    begin
      report "SIGNAL: Setting ATN to " & std_logic'image(v);
      iec_atn <= v;
    end procedure;
    procedure iec_data_out_rotate is
    begin
      -- Rotate byte being sent completely, so repeated sending
      -- of same byte is possible without having to re-write it.
      iec_data_out(6 downto 0) <= iec_data_out(7 downto 1); iec_data_out(7) <= iec_data_out(0);
    end procedure;
  begin

    if rising_edge(clock81) then
      if timing_sync_toggle /= last_timing_sync_toggle then
        last_timing_sync_toggle <= timing_sync_toggle;
        cycles <= 0;
        usecs <= 0;
      elsif cycles < (81-1) then
        cycles <= cycles + 1;
      else
        cycles <= 0;
        usec_toggle <= not usec_toggle;
        if usecs < 999 then
          usecs <= usecs + 1;
        else
          usecs <= 0;
          msec_toggle <= not msec_toggle;
        end if;
      end if;
    end if;
    
    if fastio_addr(19 downto 4) = x"d369"
      and (to_integer(fastio_addr(3 downto 0))>6)
      and (to_integer(fastio_addr(3 downto 0))<11)
      and fastio_read='1' then
      case fastio_addr(3 downto 0) is
        when x"7" => -- Read IRQ register
          fastio_rdata <= iec_irq;
        when x"8" => -- Read from status register
          fastio_rdata <= iec_status;
        when x"9" => -- Read from data register
          fastio_rdata <= iec_data;
        when x"a" => -- Read device info
          fastio_rdata <= iec_devinfo;
        when others => fastio_rdata <= (others => 'Z');
      end case;
    else
      fastio_rdata <= (others => 'Z');
    end if;
    
    if rising_edge(clock) then

      debug_state <= to_unsigned(iec_state,12);
      debug_usec <= to_unsigned(wait_usec,8);
      debug_msec <= to_unsigned(wait_msec,8);

      debug_waits(0) <= wait_clk_high;
      debug_waits(1) <= wait_clk_low;
      debug_waits(2) <= wait_data_high;
      debug_waits(3) <= wait_data_low;
      debug_waits(4) <= wait_srq_high;
      debug_waits(5) <= wait_srq_low;
      debug_waits(6) <= iec_advance;
      debug_waits(7) <= '0';
      
      -- Indicate busy status
      iec_irq(5) <= not iec_busy;
    
      -- Allow easy reading of IEC lines
      iec_status(5) <= iec_srq_i;
      iec_status(3) <= iec_clk_i;
      iec_status(2) <= iec_data_i;
      
      -- Trigger IRQ if appropriate event has occurred
      if (iec_irq(6) and iec_irq(6-4)) = '1' then
        iec_irq(7) <= '1';
      end if;
      if (iec_irq(5) and iec_irq(5-4)) = '1' then
        iec_irq(7) <= '1';
      end if;
      if (iec_irq(4) and iec_irq(4-4)) = '1' then
        iec_irq(7) <= '1';
      end if;
      if (iec_irq(7) and iec_irq(7-4)) = '1' then
        irq <= '0';
      else
        irq <= '1';
      end if;
      
      if fastio_addr(19 downto 4) = x"d369"
        and (to_integer(fastio_addr(3 downto 0))>6)
        and (to_integer(fastio_addr(3 downto 0))<11) then
        if fastio_write='1' then
          report "register write: $" & to_hexstring(fastio_wdata) & " -> reg $" & to_hexstring(fastio_addr(3 downto 0));
          case fastio_addr(3 downto 0) is
            when x"7" => -- Write to IRQ register
              -- Writing to IRQ bits clears the events
              iec_irq(7) <= iec_irq(7) and not fastio_wdata(7);
              iec_irq(6) <= iec_irq(6) and not fastio_wdata(6);
              iec_irq(5) <= iec_irq(5) and not fastio_wdata(5);
              iec_irq(4) <= iec_irq(4) and not fastio_wdata(4);
              iec_irq(3 downto 0) <= fastio_wdata(3 downto 0);
            when x"8" => -- Write to command register
              iec_cmd <= fastio_wdata;
              iec_new_cmd <= '1';
            when x"9" => -- Write to data register
              iec_data_out <= fastio_wdata;
            when x"a" => -- Write device info
            when others => null;
          end case;
        end if;
      end if;

      if iec_new_cmd='1' then
        report "IEC Command Dispatch: $" & to_hexstring(iec_cmd);
        iec_new_cmd <= '0';
        case iec_cmd is

          -- Abort existing command
          when x"00" =>
            iec_state <= 0;
            wait_clk_high <= '0'; wait_clk_low <= '0';
            wait_data_high <= '0'; wait_data_low <= '0';
            wait_srq_high <= '0'; wait_srq_low <= '0';
            wait_usec <= 0; wait_msec <= 0;
            iec_advance <= '0';
          
          -- Low-level / bitbashing commands
          when x"41" => -- ATN to +5V
            a('1');
          when x"61" => -- ATN low to 0V
            a('0');
          when x"43" => -- CLK line +5V (bitbashing)
            c('1');
          when x"63" => -- Pull CLK line low to 0V (bitbashing)
            c('0');
          when x"44" => -- DATA line to +5V (bitbashing)
            d('1');
          when x"64" => -- Pull DATA line low to 0V (bitbashing)
            d('0');
          when x"53" => -- SRQ line to +5V (bitbashing)
            s('1');
          when x"73" => -- Pull SRQ line low to 0V (bitbashing)
            s('0');
          when x"52" => -- Drive IEC reset pin 5V
            iec_reset <= '1';
          when x"72" => -- Drive IEC reset pin 0V
            iec_reset <= '0';
            

            -- Protocol level commands
          when x"30" => -- Request device attention (send data byte under attention)
            iec_dev_listening <= '1';
            iec_state <= 100;
            iec_busy <= '1';

            wait_clk_high <= '0'; wait_clk_low <= '0';
            wait_data_high <= '0'; wait_data_low <= '0';
            wait_srq_high <= '0'; wait_srq_low <= '0';
            wait_usec <= 0; wait_msec <= 0;
            iec_advance <= '0';
            
          when x"31" => -- Send byte
            iec_dev_listening <= '1';
          when x"32" => -- Receive byte
            iec_dev_listening <= '0';
          when x"33" => -- Send EOI without byte
          when x"34" => -- Send byte with EOI
          when x"35" => -- Turn around from talk to listen
            iec_dev_listening <= '0';
          when others => null;
        end case;
      end if;

      -- Update usec and msec denominated count-downs
      if usec_toggle /= last_usec_toggle then
        if wait_usec > 0 then
          report "TIME: decrementing usec counter to " & integer'image(wait_usec-1);
          wait_usec <= wait_usec - 1;
        end if;
        usec_toggle <= last_usec_toggle;
      end if;
      if msec_toggle /= last_msec_toggle then
        if wait_msec > 0 then
          report "TIME: decrementing msec counter to " & integer'image(wait_msec-1);
          wait_msec <= wait_msec - 1;
        end if;
        msec_toggle <= last_msec_toggle;
      end if;
      
      -- Advance state in IEC protocol transaction if the requirements are met
      if iec_state /= last_iec_state then
        report "iec_state = " & integer'image(iec_state)
          & ", wait_msec = " & integer'image(wait_msec)
          & ", wait_usec = " & integer'image(wait_usec)
          & ", iec_advance = " & std_logic'image(iec_advance);
        last_iec_state <= iec_state;
      end if;
      if (iec_state >0)
        and ((iec_advance='1')
             or (
               (wait_clk_low='0' or iec_clk_i='0')
               and (wait_clk_high='0' or iec_clk_i='1')
               and (wait_data_low='0' or iec_data_i='0')
               and (wait_data_high='0' or iec_data_i='1')
               and (wait_srq_low='0' or iec_srq_i='0')
               and (wait_srq_high='0' or iec_srq_i='1')
               and (wait_usec = 0)
               and (wait_msec = 0 )
               )
           )
      then
        report "Advancing to state " & integer'image(iec_state+1);
        iec_state <= iec_state + 1;
        if iec_advance='1' then
          report "iec_advance used.";
        else
          if wait_clk_high='1' then report "Used and clearing wait_clk_high"; end if;
          if wait_clk_low='1' then report "Used and clearing wait_clk_low"; end if;
          if wait_data_high='1' then report "Used and clearing wait_data_high"; end if;
          if wait_data_low='1' then report "Used and clearing wait_data_low"; end if;
          if wait_srq_high='1' then report "Used and clearing wait_srq_high"; end if;
          if wait_srq_low='1' then report "Used and clearing wait_srq_low"; end if;
          wait_clk_high <= '0'; wait_clk_low <= '0';
          wait_data_high <= '0'; wait_data_low <= '0';
          wait_srq_high <= '0'; wait_srq_low <= '0';
        end if;
        iec_advance <= '0';
      end if;
      case iec_state is
        -- IDLE state
        when 0 => null;

        -- Request attention from one or more devices
        when 100 =>

          iec_under_attention <= '0';
          
          -- DATA to 5V
          -- Ensure SRQ is released to 5V
          d('1'); s('1');

          -- Skip C= fast serial signal if a device is
          -- listening, so that it doesn't get mis-interpretted
          -- as data.
          -- XXX - Actually only required if the device supports
          -- C= fast serial?
          if iec_dev_listening='1' then
            iec_state <= 120;
          end if;

          -- Send data byte $FF using SRQ as clock to indicate our ability
          -- to do C= fast serial
        when 101 => s('1'); wait_usec <= 5;
        when 102 => s('0'); wait_usec <= 5;
        when 103 => s('1'); wait_usec <= 5;
        when 104 => s('0'); wait_usec <= 5;
        when 105 => s('1'); wait_usec <= 5;
        when 106 => s('0'); wait_usec <= 5;
        when 107 => s('1'); wait_usec <= 5;
        when 108 => s('0'); wait_usec <= 5;
        when 109 => s('1'); wait_usec <= 5;
        when 110 => s('0'); wait_usec <= 5;
        when 111 => s('1'); wait_usec <= 5;
        when 112 => s('0'); wait_usec <= 5;
        when 113 => s('1'); wait_usec <= 5;
        when 114 => s('0'); wait_usec <= 5;
        when 115 => s('1'); wait_usec <= 5;
        when 116 => s('0'); wait_usec <= 5;
          
        when 120 =>
          -- Reset all IEC lines:
          a('0'); -- ATN to 0V
          c('1'); -- CLK to 5V
          d('1'); -- DATA to 5V          
          s('1'); -- Ensure SRQ is released to 5V

          -- Clear relevant status bits
          iec_status(7) <= '0'; -- no DEVICE NOT FOUND error (yet)
          iec_status(1) <= '0'; -- No timeout
          iec_status(0) <= '0'; -- No data direction during timeout

          -- And also device info byte
          iec_devinfo(7) <= '0'; -- Device not (yet) detected
          iec_devinfo(6 downto 5) <= "00"; -- slow protocol
          -- Device ID being requested
          iec_devinfo(4 downto 0) <= iec_data_out(4 downto 0);

          -- Wait a little while before asserting CLK
          wait_usec <= 20;
          
        when 121 => 
          -- CLK to 0V
          c('0');

        when 122 =>
          -- Wait upto 1ms for DATA to go low
          wait_msec <= 1;
          report "IEC: Waiting for DATA to go low (device responding to ATN)";

        when 123 =>
          if iec_data_i = '0' then
            iec_state <= iec_state + 2; -- Proceed with ATN send
            wait_msec <= 0;
          end if;
        when 124 =>
          -- Timeout has occurred: DEVICE NOT PRESENT
          -- (actually it means that there are no devices at all)
          report "IEC: Attention timeout: No devices on bus";
          iec_state_reached <= to_unsigned(iec_state,12);
          iec_state <= 0;
          iec_devinfo <= x"00";
          iec_status(7) <= '1'; -- DEVICE NOT PRESENT
          iec_status(1) <= '1'; -- TIMEOUT OCCURRED ...
          iec_status(0) <= '1'; -- ... WHILE WE WERE TALKING          

          -- Release all IEC lines
          a('1');
          c('1');

          iec_busy <= '0';
          
        when 125 =>
          -- At least one device has responded

          c('1'); -- CLK to 5V

          -- Now wait upto 64ms for listener ready for data
          -- This period is actually unconstrained in the protcol,
          -- but we place a limit on it for now.
          wait_msec <= 64;

        when 126 =>
          if iec_data_i='1' then
            -- Listener ready for data
            iec_state <= iec_state + 2;
            wait_msec <= 0;
          end if;
        when 127 =>
          -- Timeout on listener ready for data
          
          -- Timeout has occurred: DEVICE NOT PRESENT
          -- (which is not strictly true, it's that device
          -- did not respond in time)
          iec_state_reached <= to_unsigned(iec_state,12);
          iec_state <= 0;
          iec_busy <= '0';
          iec_devinfo <= x"00";
          iec_status(7) <= '1'; -- DEVICE NOT PRESENT
          iec_status(1) <= '1'; -- TIMEOUT OCCURRED ...
          iec_status(0) <= '1'; -- ... WHILE WE WERE TALKING

          -- Release all IEC lines
          iec_atn <= '1';
          iec_clk_o <= '1'; iec_clk_en <= '1';

        when 128 =>
          -- Okay, all listeners are ready for the data byte.
          -- So send it using the slow protocol.
          -- After sending 7th bit, we do the JiffyDOS(tm) check
          -- by delaying, and waiting to see if the data line
          -- is pulled low by a device, indicating that it speaks
          -- the JiffyDOS protocol.  More on that when we get to it.

          -- Send the first 7 bits
          report "IEC: Sending data byte under ATN";
        when 129 => c('0'); d('1'); wait_usec <= 5;
        when 130 => null;
        when 131 => c('0'); d(iec_data_out(0)); wait_usec <= 15;
        when 132 => null;
        when 133 => c('1'); d(iec_data_out(0)); iec_data_out_rotate; wait_usec <= 20;
        when 134 => null;
        when 135 => c('0'); d('1'); wait_usec <= 5;
        when 136 => null;
        when 137 => c('0'); d(iec_data_out(0)); wait_usec <= 15;
        when 138 => null;
        when 139 => c('1'); d(iec_data_out(0)); iec_data_out_rotate; wait_usec <= 20;
        when 140 => null;
        when 141 => c('0'); d('1'); wait_usec <= 5;
        when 142 => null;
        when 143 => c('0'); d(iec_data_out(0)); wait_usec <= 15;
        when 144 => null;
        when 145 => c('1'); d(iec_data_out(0)); iec_data_out_rotate; wait_usec <= 20;
        when 146 => null;
        when 147 => c('0'); d('1'); wait_usec <= 5;
        when 148 => null;
        when 149 => c('0'); d(iec_data_out(0)); wait_usec <= 15;
        when 150 => null;
        when 151 => c('1'); d(iec_data_out(0)); iec_data_out_rotate; wait_usec <= 20;
        when 152 => null;
        when 153 => c('0'); d('1'); wait_usec <= 5;
        when 154 => null;
        when 155 => c('0'); d(iec_data_out(0)); wait_usec <= 15;
        when 156 => null;
        when 157 => c('1'); d(iec_data_out(0)); iec_data_out_rotate; wait_usec <= 20;
        when 158 => null;
        when 159 => c('0'); d('1'); wait_usec <= 5;
        when 160 => null;
        when 161 => c('0'); d(iec_data_out(0)); wait_usec <= 15;
        when 162 => null;
        when 163 => c('1'); d(iec_data_out(0)); iec_data_out_rotate; wait_usec <= 20;
        when 164 => null;
        when 165 => c('0'); d('1'); wait_usec <= 5;
        when 166 => null;
        when 167 => c('0'); d(iec_data_out(0)); wait_usec <= 15;
        when 168 => null;
        when 169 => c('1'); d(iec_data_out(0)); iec_data_out_rotate; wait_usec <= 20;
        when 170 => null;
           -- Now we have sent 7 bits, release data, keeping clock at 0V, and
           -- check for DATA being pulled low
        when 171 => c('0'); d('1'); wait_usec <= 500;
                    report "IEC: Performing JiffyDOS(tm) check";
        when 172 =>
          -- Data went low: device speaks JiffyDOS protocol
          if iec_data_i='0' then
            if iec_devinfo(6 downto 5) = "00" then
              report "IEC: Device supports JiffyDOS(tm) protocol. Waiting for DATA to release again.";
            end if;
            -- Record JiffyDOS capability
            iec_devinfo(6 downto 5) <= "10";
            -- Wait for DATA to be released again
            wait_usec <= 0; wait_data_high <= '1';
          end if;
        when 173 => c('0'); d(iec_data_out(0)); wait_usec <= 15;
        when 174 => null;
        when 175 => c('1'); d(iec_data_out(0)); iec_data_out_rotate; wait_usec <= 20;
        when 176 => null;
        when 177 => c('0'); d('1');
                    -- Allow device 1000usec = 1ms to acknowledge byte by
                    -- pulling data low
                    wait_msec <= 1;
                    report "IEC: Waiting for device to acknowledge byte";
        when 178 =>
          if iec_data_i='0' then
            report "IEC: Device acknowledged receipt of byte";
            iec_state <= iec_state + 2;
            wait_msec <= 0;
          end if;
        when 179 =>
          -- Timeout detected acknowledging byte

          -- Timeout has occurred: DEVICE NOT PRESENT
          -- (which is not strictly true, it's that device
          -- did not respond in time)
          report "IEC: DEVICE NOT PRESENT: Device failed to acknowledge byte";
          iec_state_reached <= to_unsigned(iec_state,12);
          iec_state <= 0;
          iec_devinfo <= x"00";
          iec_status(7) <= '1'; -- DEVICE NOT PRESENT
          iec_status(1) <= '1'; -- TIMEOUT OCCURRED ...
          iec_status(0) <= '1'; -- ... WHILE WE WERE TALKING

          iec_busy <= '0';
          
          -- Release all IEC lines
          iec_atn <= '1';
          c('1');

        when 180 =>
          -- Successfully sent byte
          report "IEC: Successfully completed sending byte under attention";
          iec_devinfo(7) <= '1';
          iec_busy <= '0';

          -- And we are still under attention
          iec_under_attention <= '1';
          iec_devinfo(4) <= '1';

          iec_state <= 0;
          
        when others => iec_state <= 0; iec_busy <= '0';
                       iec_state_reached <= to_unsigned(iec_state,12);

      end case;  
      
    end if;
  end process;
  
  
end questionable;
